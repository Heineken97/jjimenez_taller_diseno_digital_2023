module paint_VGA(
	input logic [255:0] Old_image,
	input logic [255:0] New_image,
	input logic [9:0] X, Y,
	output logic [7:0] Red, Green, Blue);
	
	logic [7:0] w_red, w_green, w_blue;
	
	//assign Red = w_red;
	//assign Blue = w_blue;
	//assign Green = w_green;
	
endmodule